--LIBRARIES
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

--ENTITY
ENTITY ARAB_COUNTER IS
	PORT (X,E,CLK,CLR,PRE:IN BIT;
      	      Q:INOUT BIT_VECTOR (1 DOWNTO 0));
END ARAB_COUNTER;

--ARCHITECTURE
ARCHITECTURE STRUCTURE OF ARAB_COUNTER IS
	
	COMPONENT ARAB_T_FF
		PORT (T, CLK, CLR, PRE : IN BIT;
		      Q:INOUT BIT);
	END COMPONENT;

SIGNAL T0,T1:BIT;

BEGIN
T0<=E;
T1<=(X XNOR Q(0)) AND (E);

A0:ARAB_T_FF PORT MAP(T0,CLK,CLR,PRE,Q(0));
A1:ARAB_T_FF PORT MAP(T1,CLK,CLR,PRE,Q(1));

END STRUCTURE;